// Forwarding Unit for pipelining CPU
module forwardUnit (
	input clk,    // Clock
	input clk_en, // Clock Enable
	input rst_n,  // Asynchronous reset active low
	
);

endmodule